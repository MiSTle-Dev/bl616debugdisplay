module DVI_CLKDIV (clkout, hclkin, resetn, calib);

output  clkout;
input  hclkin;
input  resetn;
input  calib;

CLKDIV clkdiv_inst (
    .CLKOUT(clkout),
    .HCLKIN(hclkin),
    .RESETN(resetn),
    .CALIB(calib)
);

defparam clkdiv_inst.DIV_MODE = "5";
//defparam clkdiv_inst.GSREN = "false";

endmodule
